5�d d        d    �� 
 CDflipflop�   ����2  W���                       ��  Cpin�   }����   }���0 0                  ��   �����   ����1 1                  �  ����  ����1 1                  �  W���  e���1 1                   �2  ����$  ����0 0 C2  ����        �2  }���$  }���1 1 Cp2  ����        ��   #���1  ����                       ��   �����   ����0 0                  ��   �����   ����1 1                  �  #���  ���1 1                  �  ����  ����1 1                   �1  ����#  ����0 0 B1  ���        �1  ����#  ����1 1 Bp1  ����        ��   ����2  4���                       ��   Z����   Z���0 0                  ��   r����   r���0 0                  �  ����  ����1 1                  �  4���  B���1 1                   �2  r���$  r���0 0 A2  ����        �2  Z���$  Z���1 1 Ap2  h���        ��  Cswitch#   ����/   ����9   ����l   ���� Clock    �/   ����/   ����1                    �#   ����#   ����0                     �)   ����)   ����0 0 Clock9   ����        ��  Cnand2�   �����   ����                       ��   �����   ����0 0 A�   ����        ��   �����   ����1 1 Bp�   ����         ��   �����   ����1 1                  �A   M����   )���                       �A   A���O   A���0 0 B9   O���        �A   5���O   5���1 1 Ap3   C���         ��   ;���}   ;���1 1                  �@   ����   ����                       �@   ���N   ���1 1 Cp0   ���        �@   ���N   ���1 1 Ap2   ���         ��   ���|   ���0 0                  ��   4����   ���                       ��   (����   (���1 1                  ��   ����   ���0 0                   ��   "����   "���1 1                  �F   �����   ����                       �F   ����T   ����0 0 B>   ����        �F   ����T   ����1 1 Ap8   ����         ��   �����   ����1 1                  �F   �����   l���                       �F   ����T   ����0 0 C=   ����        �F   x���T   x���1 1 Bp7   ����         ��   ~����   ~���1 1                  ��   �����   ����                       ��   �����   ����1 1                  ��   �����   ����1 1                   ��   �����   ����0 0                  �K  ���W  ����a  �����  ���� ClrAll    �K  ����K  ����1                    �W  ����W  ����0                     �Q  ���Q  ����1 0 ClrAllC  ���        ��  �����  �����  �����  ���� PreC    ��  �����  ����1 0                  ��  �����  ����0 0                   ��  �����  ����1 0 PreC�  ����        ��  8����  ,����  J����  8��� PreB    ��  ,����  ,���1                    ��  8����  8���0                     ��  2����  2���1 0 PreB�  J���        ��  �����  �����  �����  ���� PreA    ��  �����  ����1                    ��  �����  ����0                     ��  �����  ����1 0 PreA�  ����         ��  Cnet0 
 ��  Csegment)   ����)   ����L��   }����   }���L�)   �����   ����L��   �����   ����L��   Z����   Z���L�)   }����   }���L�)   ����)   }���L�)   }���)   ����L�)   Z���)   ����L��   Z���)   Z���      J�0       J�1      4   J�1  L��   �����   ����L��   �����   ����L��   �����   ����L��   �����   ����   ! J�0    # /   J�1    $ ( 0   J�1    '  	 J�1  L��   (����   ;���L��   ;����   ;���L��   ;����   ;���L��   (����   (��� +  % J�0  L��   ����   ���L��   ����   ���L��   ����   ���L��   ����   ��� ,  ) J�1  L��   �����   "���L��   "����   "���L��   "����   "���L��   �����   ����   - J�0    3   J�1  L��   �����   ����L��   �����   ����L��   �����   ����L��   �����   ���� 7  1 J�1  L��   �����   ~���L��   ~����   ~���L��   ~����   ~���L��   �����   ���� 8  5 J�0  L��   r����   ����L��   �����   ����L��   �����   ����L��   r����   r���   9 J�1  L�Q  ���Q  /���L�Q  ���Q  ���L�Q  /���  /���L�  4���  /���L�  4���  4���L�Q  ����Q  /���L�Q  ����  ����L�  ����  ����L�  ����  ����L�Q  ����Q  W���L�  W���Q  W���L�  W���  W���     = J�1  L�  ����  ����L��  ����  ����L��  �����  ����L�  ����  ����   I J�1  L�  #���  2���L��  2���  2���L��  2����  2���L�  #���  #���   E J�1  L�  ����  ����L��  �����  ����L�  ����  ����L��  ����  ����   A   jeremycastillo